library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity MatrixProcessor is
    port (
        
    );
end entity MatrixProcessor;

architecture rtl of MatrixProcessor is
    
begin
    
    
    
end architecture rtl;